module shift_right(A, S, Out);		// shift right logical module
	input [31:0] A;
	input [31:0] S;					// R[rd] = R[rt] >> shamt
	output [31:0] Out;
	wire [31:0] w1, w2, w3, w4, w5;
	
	mux2_1 m1(A[0], A[1], S[0], w1[0]);
	mux2_1 m2(A[1], A[2], S[0], w1[1]);
	mux2_1 m3(A[2], A[3], S[0], w1[2]);
	mux2_1 m4(A[3], A[4], S[0], w1[3]);
	mux2_1 m5(A[4], A[5], S[0], w1[4]);
	mux2_1 m6(A[5], A[6], S[0], w1[5]);
	mux2_1 m7(A[6], A[7], S[0], w1[6]);
	mux2_1 m8(A[7], A[8], S[0], w1[7]);
	mux2_1 m9(A[8], A[9], S[0], w1[8]);
	mux2_1 m10(A[9], A[10], S[0], w1[9]);
	mux2_1 m11(A[10], A[11], S[0], w1[10]);
	mux2_1 m12(A[11], A[12], S[0], w1[11]);
	mux2_1 m13(A[12], A[13], S[0], w1[12]);
	mux2_1 m14(A[13], A[14], S[0], w1[13]);
	mux2_1 m15(A[14], A[15], S[0], w1[14]);
	mux2_1 m16(A[15], A[16], S[0], w1[15]);
	mux2_1 m17(A[16], A[17], S[0], w1[16]);
	mux2_1 m18(A[17], A[18], S[0], w1[17]);
	mux2_1 m19(A[18], A[19], S[0], w1[18]);
	mux2_1 m20(A[19], A[20], S[0], w1[19]);
	mux2_1 m21(A[20], A[21], S[0], w1[20]);
	mux2_1 m22(A[21], A[22], S[0], w1[21]);
	mux2_1 m23(A[22], A[23], S[0], w1[22]);
	mux2_1 m24(A[23], A[24], S[0], w1[23]);
	mux2_1 m25(A[24], A[25], S[0], w1[24]);
	mux2_1 m26(A[25], A[26], S[0], w1[25]);	
	mux2_1 m27(A[26], A[27], S[0], w1[26]);
	mux2_1 m28(A[27], A[28], S[0], w1[27]);
	mux2_1 m29(A[28], A[29], S[0], w1[28]);
	mux2_1 m30(A[29], A[30], S[0], w1[29]);
	mux2_1 m31(A[30], A[31], S[0], w1[30]);
	mux2_1 m32(A[31], 1'b0, S[0], w1[31]);
	
	mux2_1 m33(w1[0], w1[2], S[1], w2[0]);
	mux2_1 m34(w1[1], w1[3], S[1], w2[1]);
	mux2_1 m35(w1[2], w1[4], S[1], w2[2]);
	mux2_1 m36(w1[3], w1[5], S[1], w2[3]);
	mux2_1 m37(w1[4], w1[6], S[1], w2[4]);
	mux2_1 m38(w1[5], w1[7], S[1], w2[5]);
	mux2_1 m39(w1[6], w1[8], S[1], w2[6]);
	mux2_1 m40(w1[7], w1[9], S[1], w2[7]);
	mux2_1 m41(w1[8], w1[10], S[1], w2[8]);
	mux2_1 m42(w1[9], w1[11], S[1], w2[9]);
	mux2_1 m43(w1[10], w1[12], S[1], w2[10]);
	mux2_1 m44(w1[11], w1[13], S[1], w2[11]);
	mux2_1 m45(w1[12], w1[14], S[1], w2[12]);
	mux2_1 m46(w1[13], w1[15], S[1], w2[13]);
	mux2_1 m47(w1[14], w1[16], S[1], w2[14]);
	mux2_1 m48(w1[15], w1[17], S[1], w2[15]);
	mux2_1 m49(w1[16], w1[18], S[1], w2[16]);
	mux2_1 m50(w1[17], w1[19], S[1], w2[17]);
	mux2_1 m51(w1[18], w1[20], S[1], w2[18]);
	mux2_1 m52(w1[19], w1[21], S[1], w2[19]);
	mux2_1 m53(w1[20], w1[22], S[1], w2[20]);
	mux2_1 m54(w1[21], w1[23], S[1], w2[21]);
	mux2_1 m55(w1[22], w1[24], S[1], w2[22]);
	mux2_1 m56(w1[23], w1[25], S[1], w2[23]);
	mux2_1 m57(w1[24], w1[26], S[1], w2[24]);
	mux2_1 m58(w1[25], w1[27], S[1], w2[25]);	
	mux2_1 m59(w1[26], w1[28], S[1], w2[26]);
	mux2_1 m60(w1[27], w1[29], S[1], w2[27]);
	mux2_1 m61(w1[28], w1[30], S[1], w2[28]);
	mux2_1 m62(w1[29], w1[31], S[1], w2[29]);
	mux2_1 m63(w1[30], 1'b0, S[1], w2[30]);
	mux2_1 m64(w1[31], 1'b0, S[1], w2[31]);

	mux2_1 m65(w2[0], w2[4], S[2], w3[0]);
	mux2_1 m66(w2[1], w2[5], S[2], w3[1]);
	mux2_1 m67(w2[2], w2[6], S[2], w3[2]);
	mux2_1 m68(w2[3], w2[7], S[2], w3[3]);
	mux2_1 m69(w2[4], w2[8], S[2], w3[4]);
	mux2_1 m70(w2[5], w2[9], S[2], w3[5]);
	mux2_1 m71(w2[6], w2[10], S[2], w3[6]);
	mux2_1 m72(w2[7], w2[11], S[2], w3[7]);
	mux2_1 m73(w2[8], w2[12], S[2], w3[8]);
	mux2_1 m74(w2[9], w2[13], S[2], w3[9]);
	mux2_1 m75(w2[10], w2[14], S[2], w3[10]);
	mux2_1 m76(w2[11], w2[15], S[2], w3[11]);
	mux2_1 m77(w2[12], w2[16], S[2], w3[12]);
	mux2_1 m78(w2[13], w2[17], S[2], w3[13]);
	mux2_1 m79(w2[14], w2[18], S[2], w3[14]);
	mux2_1 m80(w2[15], w2[19], S[2], w3[15]);
	mux2_1 m81(w2[16], w2[20], S[2], w3[16]);
	mux2_1 m82(w2[17], w2[21], S[2], w3[17]);
	mux2_1 m83(w2[18], w2[22], S[2], w3[18]);
	mux2_1 m84(w2[19], w2[23], S[2], w3[19]);
	mux2_1 m85(w2[20], w2[24], S[2], w3[20]);
	mux2_1 m86(w2[21], w2[25], S[2], w3[21]);
	mux2_1 m87(w2[22], w2[26], S[2], w3[22]);
	mux2_1 m88(w2[23], w2[27], S[2], w3[23]);
	mux2_1 m89(w2[24], w2[28], S[2], w3[24]);
	mux2_1 m90(w2[25], w2[29], S[2], w3[25]);	
	mux2_1 m91(w2[26], w2[30], S[2], w3[26]);
	mux2_1 m92(w2[27], w2[31], S[2], w3[27]);
	mux2_1 m93(w2[28], 1'b0, S[2], w3[28]);
	mux2_1 m94(w2[29], 1'b0, S[2], w3[29]);
	mux2_1 m95(w2[30], 1'b0, S[2], w3[30]);
	mux2_1 m96(w2[31], 1'b0, S[2], w3[31]);
	
	mux2_1 m97(w3[0], w3[8], S[3], w4[0]);
	mux2_1 m98(w3[1], w3[9], S[3], w4[1]);
	mux2_1 m99(w3[2], w3[10], S[3], w4[2]);
	mux2_1 m100(w3[3], w3[11], S[3], w4[3]);
	mux2_1 m101(w3[4], w3[12], S[3], w4[4]);
	mux2_1 m102(w3[5], w3[13], S[3], w4[5]);
	mux2_1 m103(w3[6], w3[14], S[3], w4[6]);
	mux2_1 m104(w3[7], w3[15], S[3], w4[7]);
	mux2_1 m105(w3[8], w3[16], S[3], w4[8]);
	mux2_1 m106(w3[9], w3[17], S[3], w4[9]);
	mux2_1 m107(w3[10], w3[18], S[3], w4[10]);
	mux2_1 m108(w3[11], w3[19], S[3], w4[11]);
	mux2_1 m109(w3[12], w3[20], S[3], w4[12]);
	mux2_1 m110(w3[13], w3[21], S[3], w4[13]);
	mux2_1 m111(w3[14], w3[22], S[3], w4[14]);
	mux2_1 m112(w3[15], w3[23], S[3], w4[15]);
	mux2_1 m113(w3[16], w3[24], S[3], w4[16]);
	mux2_1 m114(w3[17], w3[25], S[3], w4[17]);
	mux2_1 m115(w3[18], w3[26], S[3], w4[18]);
	mux2_1 m116(w3[19], w3[27], S[3], w4[19]);
	mux2_1 m117(w3[20], w3[28], S[3], w4[20]);
	mux2_1 m118(w3[21], w3[29], S[3], w4[21]);
	mux2_1 m119(w3[22], w3[30], S[3], w4[22]);
	mux2_1 m120(w3[23], w3[31], S[3], w4[23]);
	mux2_1 m121(w3[24], 1'b0, S[3], w4[24]);
	mux2_1 m122(w3[25], 1'b0, S[3], w4[25]);	
	mux2_1 m123(w3[26], 1'b0, S[3], w4[26]);
	mux2_1 m124(w3[27], 1'b0, S[3], w4[27]);
	mux2_1 m125(w3[28], 1'b0, S[3], w4[28]);
	mux2_1 m126(w3[29], 1'b0, S[3], w4[29]);
	mux2_1 m127(w3[30], 1'b0, S[3], w4[30]);
	mux2_1 m128(w3[31], 1'b0, S[3], w4[31]);
	
	mux2_1 m129(w4[0], w4[16], S[4], Out[0]);
	mux2_1 m130(w4[1], w4[17], S[4], Out[1]);
	mux2_1 m131(w4[2], w4[18], S[4], Out[2]);
	mux2_1 m132(w4[3], w4[19], S[4], Out[3]);
	mux2_1 m133(w4[4], w4[20], S[4], Out[4]);
	mux2_1 m134(w4[5], w4[21], S[4], Out[5]);
	mux2_1 m135(w4[6], w4[22], S[4], Out[6]);
	mux2_1 m136(w4[7], w4[23], S[4], Out[7]);
	mux2_1 m137(w4[8], w4[24], S[4], Out[8]);
	mux2_1 m138(w4[9], w4[25], S[4], Out[9]);
	mux2_1 m139(w4[10], w4[26], S[4], Out[10]);
	mux2_1 m140(w4[11], w4[27], S[4], Out[11]);
	mux2_1 m141(w4[12], w4[28], S[4], Out[12]);
	mux2_1 m142(w4[13], w4[29], S[4], Out[13]);
	mux2_1 m143(w4[14], w4[30], S[4], Out[14]);
	mux2_1 m144(w4[15], w4[31], S[4], Out[15]);
	mux2_1 m145(w4[16], 1'b0, S[4], Out[16]);
	mux2_1 m146(w4[17], 1'b0, S[4], Out[17]);
	mux2_1 m147(w4[18], 1'b0, S[4], Out[18]);
	mux2_1 m148(w4[19], 1'b0, S[4], Out[19]);
	mux2_1 m149(w4[20], 1'b0, S[4], Out[20]);
	mux2_1 m150(w4[21], 1'b0, S[4], Out[21]);
	mux2_1 m151(w4[22], 1'b0, S[4], Out[22]);
	mux2_1 m152(w4[23], 1'b0, S[4], Out[23]);
	mux2_1 m153(w4[24], 1'b0, S[4], Out[24]);
	mux2_1 m154(w4[25], 1'b0, S[4], Out[25]);	
	mux2_1 m155(w4[26], 1'b0, S[4], Out[26]);
	mux2_1 m156(w4[27], 1'b0, S[4], Out[27]);
	mux2_1 m157(w4[28], 1'b0, S[4], Out[28]);
	mux2_1 m158(w4[29], 1'b0, S[4], Out[29]);
	mux2_1 m159(w4[30], 1'b0, S[4], Out[30]);
	mux2_1 m160(w4[31], 1'b0, S[4], Out[31]);	
	
endmodule